

interface fadd_interface(input logic clock);

  logic reset;

  logic a,b,cin;
  logic S,Cout;

endinterface: fadd_interface